entity half_adder_1_bit is
	port(	A,B : in bit;
		S,C: out bit);
end entity;

architecture data of half_adder_1_bit is
	begin
		S <= A xor B;
		C <= A and B;
end architecture;entity half_adder_1_bit is
	port(	A,B : in bit;
		S,C: out bit);
end entity;

architecture data of half_adder_1_bit is
	begin
		S <= A xor B;
		C <= A and B;
end architecture;
